`timescale 1ns / 100ps
`default_nettype none

module top();

endmodule

`default_nettype wire
